bind sv_model blackbox_checker c0(.clk(clk), 
					  			  .rst(rst), 
								  .x(x),
								  .y(y));
						
		  
